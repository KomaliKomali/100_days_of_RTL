module NOR_2_gate_level(output Y, input A, B);
   nor(Y, A, B); 
endmodule

