module clock_buffer(input mclk,output bclk);
 
 buf b1(bclk,mclk);
 
endmodule 
  