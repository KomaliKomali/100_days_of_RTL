module data_flow(input A,B, output Y);
 assign Y = ~(A|B);
endmodule
 
 