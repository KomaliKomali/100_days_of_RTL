module NOR_gate_level(output Y, input A, B);

   nor(Y, A, B);  ////"nor" is a built-in primitive gate 
   
endmodule

